module spi_test (

);

endmodule
